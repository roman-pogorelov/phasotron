package aurora_params;

    // Aurora RX FIFO parameters
    parameter int unsigned      RX_FIFO_DEPTH   = 1024;
    parameter int unsigned      RX_FIFO_LWM     = 512;
    parameter int unsigned      RX_FIFO_HWM     = 1008;


    // Aurora TX FIFO parameters
    parameter int unsigned      TX_FIFO_DEPTH   = 1024;

endpackage: aurora_params